module tellers_to_digit
input t1 ; t2 ; t3;
output digit ; 


assign digit = t1 + t2 + t3 ;

endmodule