module sev_seg_decoder(num_in , seg);

input [3:0] num_in ;
output reg [6:0] seg ;

always @(*)
begin 
    case(num_in)
    4'h0: seg = 7'b1000000;
    4'h1: seg = 7'b1111001; 
    4'h2: seg = 7'b0100100; 
    4'h3: seg = 7'b0110000; 
    4'h4: seg = 7'b0011001; 
    4'h5: seg = 7'b0010010; 
    4'h6: seg = 7'b0000010; 
    4'h7: seg = 7'b1111000; 
    4'h8: seg = 7'b0000000; 
    4'h9: seg = 7'b0010000;   
    endcase 
end
endmodule

